module logic(
    input  wire A,
    input  wire B,
    output wire [1:0] X,
);
    wire and = A & B;
    wire or  = A | B;
    wire xor = A ^ B;

assign X = { and, xor };
endmodule
//lk;lasjdfoihqeirjtlieuyrotihgithub.o2i37rt9h3qoierutgoig2ieu4yrutgohg2o93ewup;rhkiuqyu09epujrtliu132ye0pgihliu wysedgfo;ohbwiuwe7dfu0po;bq3woi73erf70upoisb4iu5 7qwAspdhgo9wq3ueldsbfvki73u;pw.lesbndviuwpo3netg978rpbui7esujryfu7uyuj8590e4t98237y5r32y 5r2pq387y5r223i487ty53478y94578y454e3e874387545uwgr98y3i45hrpowheoir6hnkj3hporytjgk;34hyu50tpnm3kiiertgn984ikrglnhwe;ofdkhk.urewd;ofgnli8wiejrkht023qkwerltghu3wp4oekmrlkgjth4pojtlkguysrephn6iu3uy4tueoriutpowiuertpowiuertpowieurtopwieurtopiurt8903t4u3t4u9t40t43ut43ut4u03t40t43ut43u9t4309t43u093u4t09u34t09u34t093u4t0394ut093u4t093u4t09u34t0u34t09u34t093u4t09u34t09u34t09u34t09u34t09u34t093u4t09 erm what the sigma