`include "add.v"

module add8(
    input  wire [7:0] a,
    input  wire [7:0] b,
    output wire [8:0] x
);
// write your code here

endmodule
